library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_std.all;

entity paraserie is 

end paraserie;

architecture arch of paraserie is

end arch;
			