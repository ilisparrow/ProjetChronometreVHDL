library ieee;
use ieee.std_logic_1164.all;

entity structural is
end structural;

architecture arch of structural is
end arch;