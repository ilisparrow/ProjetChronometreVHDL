library ieee;
use ieee.std_logic_1164.all;

entity parite is
	port (E : in std_logic_vector (3 downto 0);
		  S : out std_logic_vector (4 downto 0));
end parite;

architecture arch1 of parite is
begin
end arch1;
