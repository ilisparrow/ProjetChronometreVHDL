library ieee;
use ieee.std_logic_1164.all;

entity compteur_tb is
end;

architecture bench of compteur_tb is



end bench;
