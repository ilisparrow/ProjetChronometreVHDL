library ieee;
use ieee.std_logic_1164.all;

entity unite_logique is
end unite_logique;

architecture arch of unite_logique is
begin
end arch;	
