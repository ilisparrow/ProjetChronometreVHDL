library ieee;
use ieee.std_logic_1164.all;

entity codeur is
end codeur;

architecture arch of codeur is
end arch;

		