library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_std.all;

entity compteur is
end compteur;

architecture arch of compteur is

end arch;