library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_std.all;

entity seriepara is 

end seriepara;

architecture arch of seriepara is

end arch;
			