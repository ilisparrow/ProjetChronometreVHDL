library ieee;
use ieee.std_logic_1164.all;

entity codeur_tb is
end;

architecture bench of codeur_tb is

end bench;