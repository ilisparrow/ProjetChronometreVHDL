library ieee;
use ieee.std_logic_1164.all;

entity compteur is
end compteur;

architecture arch of compteur is

end arch;